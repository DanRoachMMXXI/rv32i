@00000000
37 11 00 00 13 01 01 FC 23 2E 11 02 23 2C 81 02
13 04 01 04 23 26 04 FE 6F 00 80 02 03 27 C4 FE
93 07 44 FC 13 17 27 00 B3 07 F7 00 03 27 C4 FE
23 A0 E7 00 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 90 00 E3 DA E7 FC 93 07 00 00
13 85 07 00 83 20 C1 03 03 24 81 03 13 01 01 04
67 80 00 00
