`ifndef BRANCH_EVALUATOR_PKG_SV
`define BRANCH_EVALUATOR_PKG_SV

package branch_evaluator_pkg;
	`include "branch_evaluator_transaction.sv"
	`include "branch_evaluator_sequence.sv"

	`include "branch_evaluator_driver.sv"
	`include "branch_evaluator_monitor.sv"
	`include "branch_evaluator_agent.sv"
	`include "branch_evaluator_scoreboard.sv"
	`include "branch_evaluator_env.sv"
	`include "branch_evaluator_test.sv"
endpackage

`endif
