@00000000
13 01 01 FE 23 2E 11 00 23 2C 81 00 13 04 01 02
93 07 40 00 23 26 F4 FE 93 07 50 00 23 24 F4 FE
03 27 C4 FE 83 27 84 FE B3 07 F7 00 23 22 F4 FE
93 07 00 00 13 85 07 00 83 20 C1 01 03 24 81 01
13 01 01 02 67 80 00 00
