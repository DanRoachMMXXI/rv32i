`ifndef RF_WB_SELECT_PKG_SV
`define RF_WB_SELECT_PKG_SV

package rf_wb_select_pkg;
	`include "rf_wb_select_transaction.sv"
	`include "rf_wb_select_sequence.sv"

	`include "rf_wb_select_driver.sv"
	`include "rf_wb_select_monitor.sv"
	`include "rf_wb_select_agent.sv"
	`include "rf_wb_select_scoreboard.sv"
	`include "rf_wb_select_env.sv"
	`include "rf_wb_select_test.sv"
endpackage

`endif
