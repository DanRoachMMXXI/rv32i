@00000000
37 11 00 00 13 01 01 F1 23 26 11 0E 23 24 81 0E
13 04 01 0F 23 26 04 FE 6F 00 40 0B 83 27 C4 FE
13 D7 F7 41 13 77 37 00 B3 07 F7 00 93 D7 27 40
13 86 07 00 03 27 C4 FE 93 57 F7 41 93 D7 E7 01
33 07 F7 00 13 77 37 00 B3 07 F7 40 93 86 07 00
03 27 C4 FE 93 17 26 00 B3 86 D7 00 93 07 C4 F9
93 96 26 00 B3 87 F6 00 23 A0 E7 00 83 27 C4 FE
93 86 07 01 83 27 C4 FE 13 D7 F7 41 13 77 37 00
B3 07 F7 00 93 D7 27 40 13 86 07 00 03 27 C4 FE
93 57 F7 41 93 D7 E7 01 33 07 F7 00 13 77 37 00
B3 07 F7 40 13 87 07 00 93 17 26 00 33 87 E7 00
93 07 C4 F5 13 17 27 00 B3 07 F7 00 23 A0 D7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 F0 00 E3 D4 E7 F4 23 24 04 FE 6F 00 40 0D
23 22 04 FE 6F 00 40 0B 23 20 04 FE 23 2E 04 FC
6F 00 C0 06 83 27 84 FE 13 97 27 00 83 27 C4 FD
33 07 F7 00 93 07 C4 F9 13 17 27 00 B3 07 F7 00
83 A6 07 00 83 27 C4 FD 13 97 27 00 83 27 44 FE
33 07 F7 00 93 07 C4 F5 13 17 27 00 B3 07 F7 00
83 A7 07 00 93 85 07 00 13 85 06 00 EF 00 80 09
13 07 05 00 83 27 04 FE B3 87 E7 00 23 20 F4 FE
83 27 C4 FD 93 87 17 00 23 2E F4 FC 03 27 C4 FD
93 07 30 00 E3 D8 E7 F8 03 27 04 FE 83 27 84 FE
93 96 27 00 83 27 44 FE B3 86 F6 00 93 07 C4 F1
93 96 26 00 B3 87 F6 00 23 A0 E7 00 83 27 44 FE
93 87 17 00 23 22 F4 FE 03 27 44 FE 93 07 30 00
E3 D4 E7 F4 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 93 07 30 00 E3 D4 E7 F2 93 07 00 00
13 85 07 00 83 20 C1 0E 03 24 81 0E 13 01 01 0F
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 26 04 FE
6F 00 40 01 03 27 C4 FE 83 27 C4 FD B3 07 F7 00
23 26 F4 FE 83 27 84 FD 13 87 F7 FF 23 2C E4 FC
E3 92 07 FE 83 27 C4 FE 13 85 07 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00
