@00000000
37 11 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
23 2A 91 00 23 28 21 01 13 04 01 02 13 09 40 00
93 04 50 00 B3 07 99 00 23 26 F4 FE 93 07 00 00
13 85 07 00 83 20 C1 01 03 24 81 01 83 24 41 01
03 29 01 01 13 01 01 02 67 80 00 00
