module reorder_buffer #(
		parameter XLEN=32,
		// TODO: remove redundancy of TAG_WIDTH and BUF_SIZE
		// parameters, TAG_WIDTH = $clog2(BUF_SIZE).
		parameter TAG_WIDTH=8,
		parameter BUF_SIZE=64) (
	// Synchronous input signals
	input logic clk,
	input logic reset,	// active low

	// input signals for the instruciton to store in the buffer
	input logic		input_en,	// enable to read the values on the below signals
	input logic [1:0]	instruction_type_in,
	input logic [XLEN-1:0]	destination_in,
	// This interface allows a value to be stored in the ROB at the time
	// of allocation, for instructions like LUI, AUIPC, JAL, etc.
	// Since they're issued in order, nothing will be waiting for them
	//
	// Stores also may have the value immediately ready, but need to have
	// their address calculated and read from the AGU address bus.
	input logic [XLEN-1:0]	value_in,
	input logic		data_ready_in,
	input logic [XLEN-1:0]	pc_in,
	
	// common data bus signals
	input logic			cdb_valid,
	input wire [XLEN-1:0]		cdb_data,
	input wire [TAG_WIDTH-1:0]	cdb_rob_tag,
	input wire			cdb_exception,
	// branch_mispredict is a signal associated with the values on the CDB,
	// but will only be produced by branch FUs and consumed by the ROB.
	// As the name implies: has the branch being broadcast on the CDB been
	// mispredicted?  When this is stored in the ROB, it will flush all
	// subsequent instructions and update the PC to the value that
	// appeared on cdb_data (and was stored in rob_next_instruction)
	input wire			branch_mispredict,

	// memory address bus - a separate bus where the AGU sends
	// addresses to the ROB for STORES ONLY
	input logic		agu_address_valid,
	input logic [XLEN-1:0]	agu_address_data,	// the address
	input logic [XLEN-1:0]	agu_address_rob_tag,

	// flush signals - generated by the buffer_flusher (or whatever
	// I name it)
	// the flush signal is a bitmask for which each set bit clears the
	// entry at that index of the buffer
	// new_tail is the value of the new tail pointer and
	// will only be updated if |flush == 1
	// I've elected to only use these two signals to handle flushing by
	// making the assumption that flushes will only be one continuous
	// section of the buffer, from the failed instruction to the tail
	// pointer, thus only the tail pointer needs to be updated.
	input logic [BUF_SIZE-1:0]		flush,
	input logic [TAG_WIDTH-1:0]		new_tail,

	// the buffer itself
	output logic [BUF_SIZE-1:0]		rob_valid,
	output logic [BUF_SIZE-1:0][1:0]	rob_instruction_type,
	output logic [BUF_SIZE-1:0]		rob_address_valid,	// for stores only

	// destination is either the register index of rd or the memory
	// address that the value field will be written to.  whether it writes
	// to the register file or to memory is controlled by
	// instruction_type.
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_destination,
	// value stores the data that will be writted to the destination
	// field.  For ALU and memory instructions, this is the value that
	// appears on the CDB.  For branch instructions, this is PC+4, NOT the
	// value that appears on the CDB.
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_value,

	// data_ready is set either when the entry is allocated if the data is
	// already available (ex: LUI) or when the ROB tag appears on the
	// active CDB.
	output logic [BUF_SIZE-1:0]		rob_data_ready,
	output logic [BUF_SIZE-1:0]		rob_branch_mispredict,
	output logic [BUF_SIZE-1:0]		rob_exception,

	// In the event of an exception, we need to be able to update the PC
	// to whatever instruction is correct.  In the case of an exception,
	// the next instruction to be executed (thus the next value of PC) is
	// the PC of the excepting instruction.  For branches, we store the
	// correct next_instruction in this field when it appears on the CDB,
	// and update the PC if the branch was mispredicted
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_next_instruction,

	// the specific ROB entry being committed,
	// this is just rob_field[head], but I don't want to create an
	// entirely separate module to do this
	output logic		rob_commit_valid,
	output logic [1:0]	rob_commit_instruction_type,
	output logic		rob_commit_address_valid,
	output logic [XLEN-1:0]	rob_commit_destination,
	output logic [XLEN-1:0]	rob_commit_value,
	output logic		rob_commit_data_ready,
	output logic		rob_commit_branch_mispredict,
	output logic		rob_commit_exception,
	output logic [XLEN-1:0]	rob_commit_next_instruction,

	// circular buffer pointers
	// head needs to be output so that the buffer entry at head
	// can be processed when commit is set.
	// likely both head and tail will be needed for flushing the
	// buffer
	output logic [TAG_WIDTH-1:0] head,
	output logic [TAG_WIDTH-1:0] tail,

	output logic commit,
	output logic full
	);

	integer i;	// used to reset all buffer entries

	always @ (posedge clk) begin
		if (!reset) begin
			head <= 0;
			tail <= 0;

			// reset buffer contents
			// I think the only thing that matters is valid = 0
			for (i = 0; i < BUF_SIZE; i = i + 1) begin
				clear_entry(i[TAG_WIDTH-1:0]);
			end
		end else begin
			// store a new instruction in the buffer
			if (input_en) begin
				rob_valid[tail] <= 1;
				rob_instruction_type[tail] <= instruction_type_in;
				rob_destination[tail] <= destination_in;
				rob_value[tail] <= value_in;
				rob_data_ready[tail] <= data_ready_in;
				rob_next_instruction[tail] <= pc_in;

				tail <= tail + 1;
			end

			// read a value off the CDB
			if (cdb_valid && rob_valid[cdb_rob_tag]) begin
				// if an exception was broadcast on the CDB
				if (cdb_exception) begin
					// everything else is irrelevant, this
					// instrution will be flushed and retried
					rob_exception[cdb_rob_tag] <= cdb_exception;
					
					// it is critical that we do NOT
					// execute the below logic for
					// a branch because we do not want to
					// overwrite the value in
					// next_instruction since we need to
					// retry the execution of the branch.
				end
				// else if branch instruction
				else if (rob_instruction_type[cdb_rob_tag] == 'b01) begin
					// store the CDB value in
					// next_instruction (this is routed to
					// PC)
					rob_next_instruction[cdb_rob_tag] <= cdb_data;
					// check the branch_mispredict only if
					// this instruction is a branch
					rob_branch_mispredict[cdb_rob_tag] <= branch_mispredict;
				end else begin
					// else the CDB data is to be stored
					// in the register file or memory.
					rob_value[cdb_rob_tag] <= cdb_data;
				end

				rob_data_ready[cdb_rob_tag] <= 1;
			end

			// read an address off the memory address bus
			if (agu_address_valid && rob_instruction_type[agu_address_rob_tag] == 2'b11) begin
				// Load instructions use the destination field
				// of the ROB entry for the target register,
				// so we don't want to overwrite that with the
				// address to be loaded - that's stored in the
				// load buffer.
				rob_address_valid[agu_address_rob_tag] <= 1;
				rob_destination[agu_address_rob_tag] <= agu_address_data;
			end

			// instruction commit
			if (commit) begin
				clear_entry(head);
				head <= head + 1;
			end

			// clear any buffer entries specified by the flush
			// input
			for (i = 0; i < BUF_SIZE; i = i + 1) begin
				if (flush[i])
					clear_entry(i[TAG_WIDTH-1:0]);
			end

			if (|flush)
				tail <= new_tail;
		end
	end

	// if the instruction is a store, data_ready and address_valid both
	// need to be set, else just data_ready
	assign commit = rob_valid[head] && rob_data_ready[head]
					&& (rob_instruction_type[head] != 2'b11 || rob_address_valid[head] == 1);

	// the buffer is full if the entry that would be written to is already a valid entry
	assign full = rob_valid[tail];

	// values being committed if commit is set
	assign rob_commit_valid = rob_valid[head];
	assign rob_commit_instruction_type = rob_instruction_type[head];
	assign rob_commit_address_valid = rob_address_valid[head];
	assign rob_commit_destination = rob_destination[head];
	assign rob_commit_value = rob_value[head];
	assign rob_commit_data_ready = rob_data_ready[head];
	assign rob_commit_branch_mispredict = rob_branch_mispredict[head];
	assign rob_commit_exception = rob_exception[head];
	assign rob_commit_next_instruction = rob_next_instruction[head];

	function void clear_entry(logic[TAG_WIDTH-1:0] index);
		rob_valid[index] <= 0;
		rob_instruction_type[index] <= 0;
		rob_address_valid[index] <= 0;
		rob_destination[index] <= 0;
		rob_value[index] <= 0;
		rob_data_ready[index] <= 0;
		rob_branch_mispredict[index] <= 0;
		rob_exception[index] <= 0;
		rob_next_instruction[index] <= 0;
	endfunction
endmodule

// TODO: handle flushing load and store queues too
// for the load and store queues, we probably just take the ROB tags in each
// entry and subtract rob_head from them, so we can compare their age to
// rotated_oldest_exception_index to evaluate whether they need to be flushed.
// TODO: also flush reservation stations holding misspecualted instructions
// - reservation_station_reset probably takes in the flush output from this
//   module and checks if the bit at index rs_rob_tag is set
// TODO: also remember to flush instructions in the decode/RF stages
module buffer_flusher #(parameter BUF_SIZE, parameter TAG_WIDTH, parameter LDQ_SIZE, parameter STQ_SIZE) (
	// decided to not take in the valid signal for now, since I know
	// I designed the buffer to only update entries that are valid
	input logic [BUF_SIZE-1:0]	rob_branch_mispredict,
	input logic [BUF_SIZE-1:0]	rob_exception,
	input logic [TAG_WIDTH-1:0]	rob_head,
	input logic [TAG_WIDTH-1:0]	rob_tail,

	input logic [LDQ_SIZE-1:0]			ldq_valid,
	input logic [LDQ_SIZE-1:0][TAG_WIDTH-1:0]	ldq_rob_tag,
	input logic [STQ_SIZE-1:0]			stq_valid,
	input logic [STQ_SIZE-1:0][TAG_WIDTH-1:0]	stq_rob_tag,

	output logic [BUF_SIZE-1:0]	flush,
	output logic [TAG_WIDTH-1:0]	rob_new_tail,

	output logic [LDQ_SIZE-1:0]	flush_ldq,
	output logic [$clog2(LDQ_SIZE)-1:0]	ldq_new_tail,
	output logic [STQ_SIZE-1:0]	flush_stq,
	output logic [$clog2(STQ_SIZE)-1:0]	stq_new_tail
);
	// I opted to rotate both mispredicted and exception so that once the
	// index of the oldest instruction causing a flush is found, we can
	// compare it against rotated_exception to see if that instruction is
	// an exception.  This is important in determining if we need to flush
	// that instruction from the ROB.  If it's an exception, it needs to
	// be flushed from the ROB.  If it's just a branch misprediction, it
	// must remain in the ROB so that it can commit.
	logic [BUF_SIZE-1:0]	rotated_mispredict;
	logic [BUF_SIZE-1:0]	rotated_exception;
	logic [BUF_SIZE-1:0]	rotated_mispredict_or_exception;	// this is used to find the index of the ROB entry that needs to be flushed
	logic [TAG_WIDTH-1:0]	rob_rotated_tail;
	logic [BUF_SIZE-1:0]	rob_rotated_flush;

	logic			need_to_flush;	// bad name, but wasted too much time thinking of a good name
	logic [TAG_WIDTH-1:0]	rotated_oldest_exception_index;
	logic [TAG_WIDTH-1:0]	rotated_flush_start_index;	// what index does the flush actually start from?

	assign rotated_mispredict = (rob_branch_mispredict >> rob_head) | (rob_branch_mispredict << (BUF_SIZE - rob_head));
	assign rotated_exception = (rob_exception >> rob_head) | (rob_exception << (BUF_SIZE - rob_head));
	assign rotated_mispredict_or_exception = rotated_mispredict | rotated_exception;
	assign rob_rotated_tail = rob_tail - rob_head;

	lsb_priority_encoder #(.N(BUF_SIZE)) oldest_exception_finder /* idk man */ (
		.in(rotated_mispredict_or_exception),
		.out(rotated_oldest_exception_index),
		.valid(need_to_flush)
	);

	// if the instruction that caused the flush was an exception, the
	// flush begins at the index of that instruction.  if the flush was
	// caused by a branch misprediction, the flush starts at the index of
	// the instruction following the branch (the branch result is still
	// valid and thus needs to commit).
	assign rotated_flush_start_index = rotated_exception[rotated_oldest_exception_index] ? rotated_oldest_exception_index : rotated_oldest_exception_index + 1;

	integer i;
	always_comb begin
		for (i = 0; i < BUF_SIZE; i = i + 1) begin
			rob_rotated_flush[i] = (i >= rotated_flush_start_index) && (i < rob_rotated_tail)	// bound check
				&& need_to_flush;	// is there actually a need to flush
		end
	end

	assign flush = (rob_rotated_flush << rob_head) | (rob_rotated_flush >> (BUF_SIZE - rob_head));

	// the new tail is at the oldest instruction that was flushed
	assign rob_new_tail = rotated_flush_start_index + rob_head;

	// flush load queue entries
	integer ldq_index;
	always_comb begin
		for (ldq_index = 0; ldq_index < LDQ_SIZE; ldq_index = ldq_index + 1) begin
			flush_ldq[ldq_index] = (ldq_rob_tag[ldq_index] - rob_head) >= rotated_flush_start_index;
		end
		// TODO: figure out how to determine ldq_new_tail
	end

	// flush store queue entries
	integer stq_index;
	always_comb begin
		for (stq_index = 0; stq_index < STQ_SIZE; stq_index = stq_index + 1) begin
			flush_stq[stq_index] = (stq_rob_tag[stq_index] - rob_head) >= rotated_flush_start_index;
		end
		// TODO: figure out how to determine stq_new_tail
	end
	// TODO: write tests for flushing the load and store queues
endmodule
