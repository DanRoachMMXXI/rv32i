`ifndef ALU_PKG_SV
`define ALU_PKG_SV

package alu_pkg;
	`include "alu_driver.sv"
	`include "alu_transaction.sv"
endpackage

`endif
