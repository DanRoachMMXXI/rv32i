// TODO: write once src/reorder_buffer.sv is implemented
