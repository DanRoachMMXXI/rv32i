`ifndef ALU_OPERAND_SELECT_PKG_SV
`define ALU_OPERAND_SELECT_PKG_SV

package alu_operand_select_pkg;
	`include "alu_operand_select_transaction.sv"
	`include "alu_operand_select_sequence.sv"

	`include "alu_operand_select_driver.sv"
	`include "alu_operand_select_monitor.sv"
	`include "alu_operand_select_agent.sv"
	`include "alu_operand_select_scoreboard.sv"
	`include "alu_operand_select_env.sv"
	`include "alu_operand_select_test.sv"
endpackage

`endif
