`ifndef PC_SELECT_PKG_SV
`define PC_SELECT_PKG_SV

package pc_select_pkg;
	`include "pc_select_transaction.sv"
	`include "pc_select_sequence.sv"

	`include "pc_select_driver.sv"
	`include "pc_select_monitor.sv"
	`include "pc_select_agent.sv"
	`include "pc_select_scoreboard.sv"
	`include "pc_select_env.sv"
	`include "pc_select_test.sv"
endpackage

`endif
