// TODO list
// - PC update logic for predictions and executed mispredictions
module test_full_branch_fu;
	localparam XLEN = 32;
	localparam ROB_BUF_SIZE = 64;
	localparam ROB_TAG_WIDTH = $clog2(ROB_BUF_SIZE);
	localparam N_ALU_RS = 1;
	localparam N_AGU_RS = 1;
	localparam N_BRANCH_RS = 1;
	localparam TOTAL_RS = N_ALU_RS + N_AGU_RS + N_BRANCH_RS;
	localparam RAS_SIZE = 16;
	localparam LDQ_SIZE = 8;	// just need these to instantiate the buffer_flusher
	localparam STQ_SIZE = 8;

	logic clk = 0;
	logic reset = 0;

	logic [XLEN-1:0]	pc;
	logic [XLEN-1:0]	pc_plus_four;
	logic [XLEN-1:0]	pc_plus_immediate;

	// decode signals
	logic [31:0]			instruction;
	logic [XLEN-1:0]		immediate;
	control_signal_bus		control_signals_in;	// goes to route and RS

	logic	ras_push;
	logic	ras_pop;

	logic [XLEN-1:0]	ras_address_out;
	logic			ras_valid_out;

	logic [XLEN-1:0]	branch_target;

	// route signals
	logic				rs_enable;	// goes to enable of RS
	logic				stall;

	logic				rf_write_en;

	// register file outputs
	logic [XLEN-1:0]		rs1;
	logic [ROB_TAG_WIDTH-1:0]	rs1_rob_tag;
	logic				rs1_rob_tag_valid;
	logic [XLEN-1:0]		rs2;
	logic [ROB_TAG_WIDTH-1:0]	rs2_rob_tag;
	logic				rs2_rob_tag_valid;

	// reservation station input signals
	// the operands are generated by the operand_route module
	logic				q1_valid_in;
	logic [ROB_TAG_WIDTH-1:0]	q1_in;	// 0 if B_TYPE, 0 if rs1 value available, otherwise tag for rs1
	logic [XLEN-1:0]		v1_in;	// pc if B_TYPE, rs1 if JALR
	logic				q2_valid_in;
	logic [ROB_TAG_WIDTH-1:0]	q2_in;
	logic [XLEN-1:0]		v2_in;	// immediate if JALR, rs2 if B_TYPE
	logic [ROB_TAG_WIDTH-1:0]	rob_tag_in;

	// cdb arbitration
	logic [TOTAL_RS-1:0]	cdb_request;
	logic [TOTAL_RS-1:0]	cdb_permit;

	logic				rs_reset;

	logic [XLEN-1:0]		predicted_next_instruction_in;
	logic				branch_prediction_in;

	logic				cdb_valid;
	wire [XLEN-1:0]			cdb_data;
	wire [ROB_TAG_WIDTH-1:0]	cdb_rob_tag;
	wire				cdb_exception;
	wire				cdb_mispredicted;

	logic				tb_drive_cdb;	// the testbench drives the CDB, as though it were given access to do so by the CDB arbiter
	logic [XLEN-1:0]		tb_cdb_data;
	logic [ROB_TAG_WIDTH-1:0]	tb_cdb_rob_tag;

	logic [ROB_TAG_WIDTH-1:0]	q1_out;
	logic [XLEN-1:0]		v1_out;
	logic [ROB_TAG_WIDTH-1:0]	q2_out;
	logic [XLEN-1:0]		v2_out;
	control_signal_bus		control_signals_out;

	logic [XLEN-1:0]		pc_plus_four_out;
	logic [XLEN-1:0]		predicted_next_instruction_out;
	logic				branch_prediction_out;

	logic [ROB_TAG_WIDTH-1:0]	rob_tag_out;
	logic				busy;
	logic				ready_to_execute;

	logic [XLEN-1:0]		next_instruction;
	logic				redirect_mispredicted;
	logic				accept;
	logic				write_to_buffer;

	// reorder buffer inputs
	logic				alloc_rob_entry;	// generated by instruction_route

	// the reorder buffer
	logic [ROB_BUF_SIZE-1:0]		rob_valid;
	logic [ROB_BUF_SIZE-1:0][1:0]		rob_instruction_type;
	logic [ROB_BUF_SIZE-1:0]		rob_address_valid;
	logic [ROB_BUF_SIZE-1:0][XLEN-1:0]	rob_destination;
	logic [ROB_BUF_SIZE-1:0][XLEN-1:0]	rob_value;
	logic [ROB_BUF_SIZE-1:0]		rob_data_ready;
	logic [ROB_BUF_SIZE-1:0]		rob_branch_mispredict;
	logic [ROB_BUF_SIZE-1:0]		rob_exception;
	logic [ROB_BUF_SIZE-1:0][XLEN-1:0]	rob_next_instruction;

	// the instruction committing
	logic					rob_commit_valid;
	logic [1:0]				rob_commit_instruction_type;
	logic					rob_commit_address_valid;
	logic [XLEN-1:0]			rob_commit_destination;
	logic [XLEN-1:0]			rob_commit_value;
	logic					rob_commit_data_ready;
	logic					rob_commit_branch_mispredict;
	logic					rob_commit_exception;
	logic [XLEN-1:0]			rob_commit_next_instruction;

	logic [$clog2(ROB_BUF_SIZE)-1:0]	rob_head;
	logic [$clog2(ROB_BUF_SIZE)-1:0]	rob_tail;
	logic					rob_commit;
	logic					rob_full;

	logic [ROB_BUF_SIZE-1:0]		rob_flush;
	logic [$clog2(ROB_BUF_SIZE)-1:0]	rob_new_tail;

	assign cdb_data = tb_drive_cdb ? tb_cdb_data : {XLEN{1'bZ}};
	assign cdb_rob_tag = tb_drive_cdb ? tb_cdb_rob_tag : {ROB_TAG_WIDTH{1'bZ}};
	// don't think I need to drive cdb_exception or cdb_mispredicted from
	// the testbench

	assign pc_plus_four = pc + 4;
	assign pc_plus_immediate = pc + immediate;

	instruction_decode #(.XLEN(XLEN)) instruction_decode (
		.instruction(instruction),
		.immediate(immediate),
		.control_signals(control_signals_in)
	);

	// TODO: this is just temporary, need to bake this into
	// instruction_decode or something, but I'm just too over it all rn to
	// do that
	logic instruction_valid;
	always_comb begin
		case (control_signals_in.opcode)
			'b0110011,
			'b0010011,
			'b0000011,
			'b1100111,
			'b1100011,
			'b0100011,
			'b1101111,
			'b0110111,
			'b0010111:
				instruction_valid = 1;
			default:
				instruction_valid = 0;
		endcase
	end

	instruction_route #(.N_ALU_RS(N_ALU_RS), .N_AGU_RS(N_AGU_RS), .N_BRANCH_RS(N_BRANCH_RS)) route (
		.valid(instruction_valid),
		.instruction_type(control_signals_in.instruction_type),
		.ctl_alloc_rob_entry(control_signals_in.alloc_rob_entry),
		.ctl_alloc_ldq_entry(control_signals_in.alloc_ldq_entry),
		.ctl_alloc_stq_entry(control_signals_in.alloc_stq_entry),
		.rob_full(rob_full),
		.ldq_full(1'b0),
		.stq_full(1'b0),
		.flush(1'b0),	// not implemented yet
		.alu_rs_busy(1'b0),
		.agu_rs_busy(1'b0),
		.alloc_rob_entry(alloc_rob_entry),
		.alloc_ldq_entry(),
		.alloc_stq_entry(),
		.branch_rs_busy(busy),
		.alu_rs_route(),
		.agu_rs_route(),
		.branch_rs_route(rs_enable),
		.stall(stall)
	);

	operand_route #(.XLEN(XLEN), .ROB_SIZE(ROB_BUF_SIZE), .ROB_TAG_WIDTH(ROB_TAG_WIDTH)) operand_route (
		.opcode(control_signals_in.opcode),
		.rs1(rs1),
		.rs1_rob_tag(rs1_rob_tag),
		.rs1_rob_tag_valid(rs1_rob_tag_valid),
		.rs2(rs2),
		.rs2_rob_tag(rs2_rob_tag),
		.rs2_rob_tag_valid(rs2_rob_tag_valid),
		.pc(pc),
		.immediate(immediate),
		.rob_value(rob_value),
		.rob_data_ready(rob_data_ready),
		.q1_valid(q1_valid_in),
		.q1(q1_in),
		.v1(v1_in),
		.q2_valid(q2_valid_in),
		.q2(q2_in),
		.v2(v2_in)
	);

	cdb_arbiter #(.N(N_ALU_RS + N_AGU_RS + N_BRANCH_RS)) cdb_arbiter (
		.request(cdb_request),
		.grant(cdb_permit),
		.cdb_valid(cdb_valid)
	);

	register_file #(.XLEN(XLEN), .ROB_TAG_WIDTH(ROB_TAG_WIDTH)) rf (
		.clk(clk),
		.reset(reset),
		.rs1_index(control_signals_in.rs1_index),
		.rs2_index(control_signals_in.rs2_index),
		.alloc_rob_entry(alloc_rob_entry),
		.rob_alloc_rd_index(control_signals_in.rd_index),
		.rob_alloc_tag(rob_tail),
		.rd_index(rob_commit_destination[4:0]),
		.rd(rob_commit_value),
		.rd_rob_index(rob_head),
		.write_en(rf_write_en),
		.rs1(rs1),
		.rs1_rob_tag(rs1_rob_tag),
		.rs1_rob_tag_valid(rs1_rob_tag_valid),
		.rs2(rs2),
		.rs2_rob_tag(rs2_rob_tag),
		.rs2_rob_tag_valid(rs2_rob_tag_valid)
	);

	ras_control ras_control (
		.jump(control_signals_in.jump),
		.jalr(control_signals_in.jalr),
		.rs1_index(control_signals_in.rs1_index),
		.rd_index(control_signals_in.rd_index),

		.push(ras_push),
		.pop(ras_pop)
	);

	return_address_stack #(.XLEN(XLEN), .STACK_SIZE(RAS_SIZE)) ras (
		.clk(clk),
		.reset(reset),

		.address_in(pc_plus_four),
		.push(ras_push),
		.pop(ras_pop),

		// not doing checkpointing in this test yet, as it's already
		// covered in the unit test
		.checkpoint(),
		.restore_checkpoint(),

		.address_out(ras_address_out),
		.valid_out(ras_valid_out),

		// debug signals, no need to attach these unless shit hits the
		// fan
		.stack(),
		.stack_valid(),
		.stack_pointer(),
		.sp_checkpoint()
	);

	branch_target #(.XLEN(XLEN)) branch_target_calculator (
		.pc(pc),
		// TODO: for now, I'm assuming that we only use the values on
		// the RAS to predict values for JALR instructions.  as noted
		// in cpu.sv, I may cache or forward values from LUI and AUIPC
		// if the registers match. If I do, I should update this test.
		// Until then, JALR predictions that don't pop off the stack
		// will use 0 as the source, which is just as useless as any
		// other number, but for the purposes of testing the branch
		// pipeline I'm down with it as it is near guaranteed to
		// mispredict and I can validate that it flushes.
		.rs1(ras_address_out),
		.immediate(immediate),
		.jalr(control_signals_in.jalr),

		.branch_target(branch_target)
	);

	branch_predictor #(.XLEN(XLEN)) branch_predictor (
		.pc_plus_four(pc_plus_four),
		.branch_target(branch_target),
		.jump(control_signals_in.jump),
		.branch(control_signals_in.branch),
		.branch_predicted_taken(branch_prediction_in)
	);

	reservation_station #(.XLEN(XLEN), .TAG_WIDTH(ROB_TAG_WIDTH)) reservation_station (
		.clk(clk),
		.reset(rs_reset),
		.enable(rs_enable),
		.dispatched_in(accept),
		.q1_valid_in(q1_valid_in),
		.q1_in(q1_in),
		.v1_in(v1_in),
		.q2_valid_in(q2_valid_in),
		.q2_in(q2_in),
		.v2_in(v2_in),
		.control_signals_in(control_signals_in),
		.rob_tag_in(rob_tag_in),	// this needs to get rob.write_to routed to it somehow
		.pc_plus_four_in(pc_plus_four),
		.predicted_next_instruction_in(predicted_next_instruction_in),
		.branch_prediction_in(branch_prediction_in),
		.cdb_valid(cdb_valid),
		.cdb_rob_tag(cdb_rob_tag),
		.cdb_data(cdb_data),
		.q1_valid_out(),
		.q1_out(q1_out),
		.v1_out(v1_out),
		.q2_valid_out(),
		.q2_out(q2_out),
		.v2_out(v2_out),
		.control_signals_out(control_signals_out),
		.rob_tag_out(rob_tag_out),
		.pc_plus_four_out(pc_plus_four_out),
		.predicted_next_instruction_out(predicted_next_instruction_out),
		.branch_prediction_out(branch_prediction_out),
		.busy(busy),
		.ready_to_execute(ready_to_execute)
	);

	reservation_station_reset #(.TAG_WIDTH(ROB_TAG_WIDTH)) reservation_station_reset (
		.global_reset(reset),
		.bus_valid(cdb_valid),
		.bus_rob_tag(cdb_rob_tag),
		.rs_rob_tag(rob_tag_out),
		.reservation_station_reset(rs_reset)
	);

	branch_functional_unit #(.XLEN(XLEN)) fu (
		.v1(v1_out),
		.v2(v2_out),
		.pc_plus_four(pc_plus_four_out),
		.pc_plus_immediate(pc_plus_immediate),
		.predicted_next_instruction(predicted_next_instruction_out),
		.funct3(control_signals_out.funct3),
		.jalr(control_signals_out.jalr),
		.branch(control_signals_out.branch),
		.next_instruction(next_instruction),
		.redirect_mispredicted(redirect_mispredicted),
		.ready_to_execute(ready_to_execute),
		.accept(accept),
		.write_to_buffer(write_to_buffer)
	);

	functional_unit_output_buffer #(.XLEN(XLEN), .TAG_WIDTH(ROB_TAG_WIDTH)) output_buf (
		.clk(clk),
		.reset(reset),
		.value(next_instruction),
		.tag(rob_tag_out),
		.exception(1'b0),	// TODO: actually do something with this
		.redirect_mispredicted(redirect_mispredicted),
		.write_en(write_to_buffer),
		.not_empty(cdb_request[0]),
		.data_bus_permit(cdb_permit[0]),
		.data_bus_data(cdb_data),
		.data_bus_tag(cdb_rob_tag),
		.data_bus_exception(cdb_exception),
		.data_bus_redirect_mispredicted(cdb_mispredicted),
		.read_from(),
		.write_to()
	);

	reorder_buffer #(.XLEN(XLEN), .TAG_WIDTH(ROB_TAG_WIDTH), .BUF_SIZE(ROB_BUF_SIZE)) rob (
		.clk(clk),
		.reset(reset),
		.input_en(alloc_rob_entry),
		.instruction_type_in(control_signals_in.instruction_type),
		// TODO: these signals
		.destination_in(),
		.value_in(),
		.data_ready_in(),
		.pc_in(pc),
		.cdb_valid(cdb_valid),
		.cdb_data(cdb_data),
		.cdb_rob_tag(cdb_rob_tag),
		.cdb_exception(cdb_exception),
		.branch_mispredict(cdb_mispredicted),
		.agu_address_valid(),
		.agu_address_data(),
		.agu_address_rob_tag(),
		.flush(rob_flush),
		.new_tail(rob_new_tail),
		.rob_valid(rob_valid),
		.rob_instruction_type(rob_instruction_type),
		.rob_address_valid(rob_address_valid),
		.rob_destination(rob_destination),
		.rob_value(rob_value),
		.rob_data_ready(rob_data_ready),
		.rob_branch_mispredict(rob_branch_mispredict),
		.rob_exception(rob_exception),
		.rob_next_instruction(rob_next_instruction),
		.rob_commit_valid(rob_commit_valid),
		.rob_commit_instruction_type(rob_commit_instruction_type),
		.rob_commit_address_valid(rob_commit_address_valid),
		.rob_commit_destination(rob_commit_destination),
		.rob_commit_value(rob_commit_value),
		.rob_commit_data_ready(rob_commit_data_ready),
		.rob_commit_branch_mispredict(rob_commit_branch_mispredict),
		.rob_commit_exception(rob_commit_exception),
		.rob_commit_next_instruction(rob_commit_next_instruction),
		.head(rob_head),
		.tail(rob_tail),
		.commit(rob_commit),
		.full(rob_full)
	);

	buffer_flusher #(.BUF_SIZE(ROB_BUF_SIZE), .TAG_WIDTH(ROB_TAG_WIDTH), .LDQ_SIZE(LDQ_SIZE), .STQ_SIZE(STQ_SIZE)) buffa_flusha (
		.rob_branch_mispredict(rob_branch_mispredict),
		.rob_exception(rob_exception),
		.rob_head(rob_head),
		.rob_tail(rob_tail),

		// at the time of writing this test these don't even do
		// anything, and will probably change once I implement the
		// flushing of the load and store queues
		.ldq_valid(),
		.ldq_rob_tag(),
		.stq_valid(),
		.stq_rob_tag(),

		.flush(rob_flush),
		.rob_new_tail(rob_new_tail),

		.flush_ldq(),
		.ldq_new_tail(),
		.flush_stq(),
		.stq_new_tail()
	);

	rf_writeback rf_writeback (
		.rob_commit(rob_commit),
		.rob_commit_valid(rob_commit_valid),
		.rob_commit_instruction_type(rob_commit_instruction_type),
		.rob_commit_exception(rob_commit_exception),
		.rf_write_en(rf_write_en)
	);

	// disable the active low reset after the first clock cycle
	initial begin
		#10 reset = 1;
	end

	always begin
		#5 clk = ~clk;
	end

	initial begin	// test logic
		# 10	// wait for reset

		// TODO: eventually, this is going to break, as I don't intend
		// to execute JAL in the FU.  It will automatically just jump
		// to the computed PC
		pc = 'hC;
		instruction = 'h0140006f;	// jal x0, 20
		# 2
		assert(immediate == 20);
		assert(ras_push == 0);
		assert(ras_pop == 0);
		assert(ras_valid_out == 0);
		assert(branch_target == 'hC + 20);

		# 8
		assert(ready_to_execute == 1);
		assert(busy == 1);
		assert(stall == 1);	// we never changed instruction, so it would be trying to issue it again
		assert(write_to_buffer == 1);
		# 10
		assert(cdb_request == 'b1);
		assert(cdb_permit == 'b1);
		assert(cdb_valid == 1);
		// cdb_data is 0 because no logic in the FU actually handles JAL
		assert(busy == 1);	// on the next cycle, the RS will see its ROB tag on the CDB and clear itself
		# 10

		// instruction = 'h00000013;	// addi x0, x0, 0 - conventional NOP
		instruction = 0;	// cleared instruction - unconventional NOP, but must do nothing
		assert(busy == 0);
		assert(rob_valid[0] == 'b1);
		assert(rob_commit == 1);
		assert(rf_write_en == 1);	// doesn't really matter if this is set or clear, rd = x0 and won't be updated in the RF

		# 10
		assert(rob_valid == 0);
		assert(rob_commit == 0);

		// instruction = 'hFEDFF06F;	// jal x0, -20
		# 10
		$display("All assertions passed.");
		$finish();
	end
endmodule
