typedef struct packed {
	logic branch_predicted_taken;
	logic branch_mispredicted;
} branch_signal_bus;
