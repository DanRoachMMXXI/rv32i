/*
 * TODO: be mentally prepared to handle flushing mispredicts
 * it might not be too bad if done simply: flush all instructions when the
 * branch result commits.  that would be very inefficient tho, because we want
 * to flush and start fetching new instructions as soon as we know the branch
 * was incorrect.  We can't use the pc value to determine if an instruciton
 * was executed on a misprediction.  We need to leverage the ordering of
 * instructions in the buffer.  So for all elements after the mispredicted
 * branch (and before the head index), they need to be flushed.
 * [ valid, tail, empty, empty, head, valid, mispredicted, valid ]
 *     0       1        2      3        4        5         6          7
 * in this example, indices 7 and 0 would need to be flushed when we find out
 * that the branch prediction was wrong.  reminder that 1 is not yet occupied.
 * we can guarantee that a mispredicted instruciton is between head and
 * tail, but I don't know if that guarantee is useful in implementing the
 * logic.
 *
 * we can not guarantee that mispredicted != tail.  they are equal if the
 * buffer is full and the mispredicted branch is the first in the buffer, and
 * every other instruction in the buffer is flushed.
 *
 * the instructions to flush are the instructions between the index of the
 * mispredicted index and the tail index, not inclusive.
 * 
 * The textbook DOES say that the buffer flushing is done when the
 * mispredicted branch commits.  I think my assessment is still correct, but
 * it may be a good idea to implement the simple and suboptimal solution
 * quickly to get it done, then fuck about with more complicated
 * optimizations.
 * The textbook then ALSO does say in practice processors do what I described
 * above.  Plan is probably still valid: do easy thing, then hard thing.
 *
 * It may become easier to offload the flushing of the buffer to another
 * component, and take in the signals to flush specific entries of the buffer.
 */
module reorder_buffer #(
		parameter XLEN=32,
		// TODO: remove redundancy of TAG_WIDTH and BUF_SIZE
		// parameters, TAG_WIDTH = $clog2(BUF_SIZE).
		parameter TAG_WIDTH=8,
		parameter BUF_SIZE=64) (
	// Synchronous input signals
	input logic clk,
	input logic reset,	// active low

	// input signals for the instruciton to store in the buffer
	input logic		input_en,	// enable to read the values on the below signals
	input logic [1:0]	instruction_type_in,
	input logic [XLEN-1:0]	destination_in,
	// This interface allows a value to be stored in the ROB at the time
	// of allocation, for instructions like LUI, AUIPC, JAL, etc.
	// Since they're issued in order, nothing will be waiting for them
	//
	// Stores also may have the value immediately ready, but need to have
	// their address calculated and read from the AGU address bus.
	input logic [XLEN-1:0]	value_in,
	input logic		data_ready_in,
	input logic [XLEN-1:0]	next_instruction_in,
	
	// common data bus signals
	input logic			cdb_valid,
	input wire [XLEN-1:0]		cdb_data,
	input wire [TAG_WIDTH-1:0]	cdb_rob_tag,
	input wire			cdb_exception,

	// memory address bus - a separate bus where the AGU sends
	// addresses to the ROB for STORES ONLY
	input logic		agu_address_valid,
	input logic [XLEN-1:0]	agu_address_data,	// the address
	input logic [XLEN-1:0]	agu_address_rob_tag,

	// flush signals - generated by the rob_exception_handler (or whatever
	// I name it)
	// the flush signal is a bitmask for which each set bit clears the
	// entry at that index of the buffer
	// new_tail is the value of the new tail pointer and
	// will only be updated if |flush == 1
	// I've elected to only use these two signals to handle flushing by
	// making the assumption that flushes will only be one continuous
	// section of the buffer, from the failed instruction to the tail
	// pointer, thus only the tail pointer needs to be updated.
	input logic [BUF_SIZE-1:0]		flush,
	input logic [TAG_WIDTH-1:0]		new_tail,

	// the buffer itself
	output logic [BUF_SIZE-1:0]		rob_valid,
	output logic [BUF_SIZE-1:0][1:0]	rob_instruction_type,
	output logic [BUF_SIZE-1:0]		rob_address_valid,	// for stores only

	// destination is either the register index of rd or the memory
	// address that the value field will be written to.  whether it writes
	// to the register file or to memory is controlled by
	// instruction_type.
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_destination,
	// value stores the data that will be writted to the destination
	// field.  For ALU and memory instructions, this is the value that
	// appears on the CDB.  For branch instructions, this is PC+4, NOT the
	// value that appears on the CDB.
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_value,

	// data_ready is set either when the entry is allocated if the data is
	// already available (ex: LUI) or when the ROB tag appears on the
	// active CDB.
	output logic [BUF_SIZE-1:0]		rob_data_ready,
	output logic [BUF_SIZE-1:0]		rob_exception,

	// In the event of an exception, we need to be able to restore the PC
	// to the correct next instruction.  For ALU/memory instructions, this
	// is just pc_plus_four.  For branches, if there's a mispredict, we
	// store the correct next_instruction in here and update PC like any
	// other exception.
	output logic [BUF_SIZE-1:0][XLEN-1:0]	rob_next_instruction,

	// circular buffer pointers
	// head needs to be output so that the buffer entry at head
	// can be processed when commit is set.
	// likely both head and tail will be needed for flushing the
	// buffer
	output logic [TAG_WIDTH-1:0] head,
	output logic [TAG_WIDTH-1:0] tail,

	output logic commit,
	output logic full
	);

	integer i;	// used to reset all buffer entries

	always @ (posedge clk) begin
		if (!reset) begin
			head <= 0;
			tail <= 0;

			// reset buffer contents
			// I think the only thing that matters is valid = 0
			for (i = 0; i < BUF_SIZE; i = i + 1) begin
				clear_entry(i[TAG_WIDTH-1:0]);
			end
		end else begin
			// store a new instruction in the buffer
			if (input_en) begin
				rob_valid[tail] <= 1;
				rob_instruction_type[tail] <= instruction_type_in;
				rob_destination[tail] <= destination_in;
				rob_value[tail] <= value_in;
				rob_data_ready[tail] <= data_ready_in;

				tail <= tail + 1;
			end

			// read a value off the CDB
			if (cdb_valid && rob_valid[cdb_rob_tag]) begin
				// if branch instruction
				if (rob_instruction_type[cdb_rob_tag] == 'b01) begin
					// store the CDB value in
					// next_instruction (this is routed to
					// PC)
					rob_next_instruction[cdb_rob_tag] <= cdb_data;
				end else begin
					// else the CDB data is to be stored
					// in the register file or memory.
					rob_value[cdb_rob_tag] <= cdb_data;
				end

				rob_data_ready[cdb_rob_tag] <= 1;
				rob_exception[cdb_rob_tag] <= cdb_exception;
			end

			// read an address off the memory address bus
			if (agu_address_valid && rob_instruction_type[agu_address_rob_tag] == 2'b11) begin
				// Load instructions use the destination field
				// of the ROB entry for the target register,
				// so we don't want to overwrite that with the
				// address to be loaded - that's stored in the
				// load buffer.
				rob_address_valid[agu_address_rob_tag] <= 1;
				rob_destination[agu_address_rob_tag] <= agu_address_data;
			end

			// instruction commit
			if (commit) begin
				clear_entry(head);
				head <= head + 1;
			end

			// clear any buffer entries specified by the flush
			// input
			for (i = 0; i < BUF_SIZE; i = i + 1) begin
				if (flush[i])
					clear_entry(i[TAG_WIDTH-1:0]);
			end

			if (|flush)
				tail <= new_tail;
		end
	end

	// if the instruction is a store, data_ready and address_valid both
	// need to be set, else just data_ready
	assign commit = rob_valid[head] && rob_data_ready[head]
					&& (rob_instruction_type[head] != 2'b11 || rob_address_valid[head] == 1);

	// the buffer is full if the entry that would be written to is already a valid entry
	assign full = rob_valid[tail];

	function void clear_entry(logic[TAG_WIDTH-1:0] index);
		rob_valid[index] <= 0;
		rob_instruction_type[index] <= 0;
		rob_address_valid[index] <= 0;
		rob_destination[index] <= 0;
		rob_value[index] <= 0;
		rob_data_ready[index] <= 0;
		rob_exception[index] <= 0;
		rob_next_instruction[index] <= 0;
	endfunction
endmodule

// TODO: I'm probably misusing the phrase "exception".  Page 20 of the RISC-V
// Unprivileged ISA gives some clarity into what exceptions are and how
// they're handled.  Branch misprediction and order failures do not seem to
// fall into the category of exceptions
// "The general behavior of most RISC-V EEIs is that a trap to some handler
// occurs when an exception is signaled on an instruction"
// I suppose we shall refer to these as misspeculations?  something
// branch mispredictions: we DO want to commit these instructions
// load ordering failures: we do NOT want to commit these, we need to retry
// the instruction before it can be committed
// BOOM says it treats ordering failures as exceptions, but it only causes
// a pipeline retry
// The Load/Store unit can incur two exceptions:
// - page faults
// - load ordering failures
// while I am not using virtual memory (yet), I assume these both yield the
// same result: retry the operation.
// The Branch unit can incur one exception: misalignment
// I guess everything that is an exception gets retried in the pipeline (how
// tf do I do that?).  Branch mispreidction just flushes everything after it,
// no retry tho.
//
// TODO: handle flushing load and store queues too
// for the load and store queues, we probably just take the ROB tags in each
// entry and subtract rob_head from them, so we can compare their age to
// rotated_oldest_exception_index to evaluate whether they need to be flushed.
//
// I THINK I AM GOING TO KEEP THIS MODULE RELATED TO FLUSHING THE ROB, NOT
// HANDLING EXCEPTIONS, SO TODO RENAME THIS MODULE rob_flush_generator OR
// SOMETHING
module rob_exception_handler #(parameter BUF_SIZE, parameter TAG_WIDTH) (
	// decided to not take in the valid signal for now, since I know
	// I designed the buffer to only update entries that are valid
	input logic [BUF_SIZE-1:0]	rob_exception,
	input logic [TAG_WIDTH-1:0]	rob_head,
	input logic [TAG_WIDTH-1:0]	rob_tail,
	// TODO: inputs from LDQ and STQ

	output logic [BUF_SIZE-1:0]	flush,
	output logic [TAG_WIDTH-1:0]	new_tail
	// output logic [LDQ_SIZE-1:0]	flush_ldq,
	// output logic [$clog2(LDQ_SIZE)-1:0]	ldq_new_tail,
	// output logic [STQ_SIZE-1:0]	flush_stq,
	// output logic [$clog2(STQ_SIZE)-1:0]	stq_new_tail
);
	logic [BUF_SIZE-1:0]	rob_rotated_exception;
	logic [TAG_WIDTH-1:0]	rob_rotated_tail;
	logic [BUF_SIZE-1:0]	rob_rotated_flush;

	logic			exception;
	logic [TAG_WIDTH-1:0]	rotated_oldest_exception_index;

	assign rob_rotated_exception = (rob_exception >> rob_head) | (rob_exception << (BUF_SIZE - rob_head));
	assign rob_rotated_tail = rob_tail - rob_head;

	lsb_priority_encoder #(.N(BUF_SIZE)) oldest_exception_finder /* idk man */ (
		.in(rob_rotated_exception),
		.out(rotated_oldest_exception_index),
		.valid(exception)
	);

	integer i;
	always_comb begin
		for (i = 0; i < BUF_SIZE; i = i + 1) begin
			// flush entries that are between the index of the
			// oldest exception index (exclusive?) and the tail
			// (exclusive) ONLY IF there is actually an exception
			// (indicated by the exception signal)
			rob_rotated_flush[i] = (i > rotated_oldest_exception_index) && (i < rob_rotated_tail) && exception;
		end
	end

	assign flush = (rob_rotated_flush << rob_head) | (rob_rotated_flush >> (BUF_SIZE - rob_head));
endmodule
