/*
 * Tracks in flight load operations
 * so wtf does this thing need to do:
 * - allocate entries new load instructions (DONE)
 *   - set valid bit (DONE)
 *   - probably store ROB tag as an identifier? (DONE)
 * - store addresses from AGU
 *   - update entry with address and set address_valid (DONE)
 *   - fire load as soon as address arrives
 * - update load entries
 *   - mark loads as sent
 *   - cancel loads with dependent stores
 *   - update all the other signals in load_queue_entry
 * - compare against store addresses once address arrives
 *   - THIS IS ALL DONE WITH A SEPARATE COMPONENT
 *   - if there's a match
 *	- cancel the fired load operation
 *	- forward the data if it's available in the store buffer
 *	- sleep until the data is available if it isn't already available
 */
module load_queue 
	import lsu_pkg::*;
	/* #(parameter XLEN=32, parameter ROB_TAG_WIDTH=32, parameter LDQ_SIZE=16, parameter STQ_SIZE=16) */ (
	input logic clk,
	input logic reset,

	// signals to allocate a new load instruction
	// tentatively planning to use the ROB tag to track incoming updates
	// to this load.
	// - address from the AGU
	// - load completed from memory (tracked by caches)
	// also thinking I need the ROB tag to broadcast to the CDB, but
	// I need to figure out what component is responsible for broadcasting
	input logic alloc_ldq_entry,
	input logic [ROB_TAG_WIDTH-1:0] rob_tag_in,

	// signals to store addresses from an AGU
	input logic agu_address_valid,
	input logic [XLEN-1:0] agu_address_data,
	input logic [ROB_TAG_WIDTH-1:0] agu_address_rob_tag,	// use to identify which

	// signals to indicate a load has been fired
	input logic load_executed,
	input logic [ROB_TAG_WIDTH-1:0] load_executed_rob_tag,

	// signals from the memory interface to designate a succeeded load
	// the load_succeeded_rob_tag is tracked by cache miss registers in
	// the caches
	input logic load_succeeded,				// bool to say if a load succeeded
	input logic [ROB_TAG_WIDTH-1:0] load_succeeded_rob_tag,	// ROB tag of the succeeded load

	input logic set_store_mask,	// bool to set a store mask
	input logic [STQ_SIZE-1:0] store_mask,
	input logic [$clog2(LDQ_SIZE)-1:0] store_mask_index,	// TODO might be ROB tag idk

	// rob signals to know when loads commit
	// loads are stored in program order so we know we're freeing the head
	input logic rob_commit,
	input logic rob_commit_type,

	input logic set_order_fail,	// signals that an order failure was detected
	input logic [$clog2(LDQ_SIZE)-1:0] order_fail_index,	// LDQ index of the load that experienced the order failure

	output load_queue_entry [LDQ_SIZE-1:0] load_queue_entries
	);

	// circular buffer pointers
	logic [$clog2(LDQ_SIZE)-1:0] head;
	logic [$clog2(LDQ_SIZE)-1:0] tail;

	integer i;

	always_ff @ (posedge clk) begin
		if (!reset) begin
			head <= 0;
			tail <= 0;

			for (i = 0; i < LDQ_SIZE; i = i + 1) begin
				clear_entry(i);
			end
		end else begin
			// place a new load instruction in the load buffer
			if (alloc_ldq_entry) begin
				load_queue_entries[tail].valid <= 1;
				load_queue_entries[tail].rob_tag <= rob_tag_in;
				tail <= tail + 1;
			end

			// set order failure if it was detected by the searcher
			if (set_order_fail) begin
				load_queue_entries[order_fail_index].order_fail <= 1;
			end

			// set the store mask generated by the searcher at the specified index
			if (set_store_mask) begin
				load_queue_entries[store_mask_index].store_mask <= store_mask;
			end

			// if the ROB committed a load, free the load at the head
			if (rob_commit && rob_commit_type == 0) begin
				clear_entry(head);
				head <= head + 1;
			end

			// TODO:
			// - order_fail
			//	- "To discover ordering failures, when a store
			//	commits, it checks the entire LDQ for any
			//	address matches. If there is a match, the
			//	store checks to see if the load has executed,
			//	and if it got its data from memory or if the
			//	data was forwarded from an older store. In
			//	either case, a memory ordering failure has
			//	occurred."
			//	- needs to be able to update all or multiple
			//	entries in one cycle
			// - forward_stq_data
			// - forward_stq_index

			// loop to do operations on every entry
			for (i = 0; i < LDQ_SIZE; i = i + 1) begin	// each entry in the buffer makes this comparison
				// READ ADDRESS FROM THE AGU
				// if the address from the AGU is to be read and the ROB tag matches
				if (load_queue_entries[i].valid && agu_address_valid && agu_address_rob_tag == load_queue_entries[i].rob_tag) begin
					// if match, update address and declare it to be valid
					load_queue_entries[i].address <= agu_address_data;
					load_queue_entries[i].address_valid <= 1;
				end

				if (load_queue_entries[i].valid && load_executed && load_executed_rob_tag == load_queue_entries[i].rob_tag) begin
					load_queue_entries[i].executed <= 1;
				end

				if (load_queue_entries[i].valid && load_succeeded && load_succeeded_rob_tag == load_queue_entries[i].rob_tag) begin
					load_queue_entries[i].succeeded <= 1;
				end
			end
		end
	end

	function clear_entry(logic[$clog2(LDQ_SIZE)-1:0] index);
		load_queue_entries[index].valid <= 0;
		load_queue_entries[index].address <= 0;
		load_queue_entries[index].address_valid <= 0;
		load_queue_entries[index].executed <= 0;
		load_queue_entries[index].succeeded <= 0;
		load_queue_entries[index].order_fail <= 0;
		load_queue_entries[index].store_mask <= 0;
		load_queue_entries[index].forward_stq_data <= 0;
		load_queue_entries[index].forward_stq_index <= 0;
		load_queue_entries[index].rob_tag <= 0;
	endfunction
endmodule
