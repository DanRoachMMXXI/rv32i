/*
 * Tracks in flight load operations
 * so wtf does this thing need to do:
 * - allocate entries new load instructions (DONE)
 *   - set valid bit (DONE)
 *   - probably store ROB tag as an identifier? (DONE)
 * - store addresses from AGU
 *   - update entry with address and set address_valid (DONE)
 *   - fire load as soon as address arrives
 * - update load entries
 *   - mark loads as sent
 *   - cancel loads with dependent stores
 *   - update all the other signals in load_queue_entry
 * - compare against store addresses once address arrives
 *   - THIS IS ALL DONE WITH A SEPARATE COMPONENT
 *   - if there's a match
 *	- cancel the fired load operation
 *	- forward the data if it's available in the store buffer
 *	- sleep until the data is available if it isn't already available
 */
module load_queue 
	import lsu_pkg::*;
	/* #(parameter XLEN=32, parameter ROB_TAG_WIDTH=32, parameter LDQ_SIZE=16, parameter STQ_SIZE=16) */ (
	input logic clk,
	input logic reset,

	// signals to allocate a new load instruction
	// tentatively planning to use the ROB tag to track incoming updates
	// to this load.
	// - address from the AGU
	// - load completed from memory (tracked by caches)
	// also thinking I need the ROB tag to broadcast to the CDB, but
	// I need to figure out what component is responsible for broadcasting
	input logic alloc_ldq_entry,
	input logic [ROB_TAG_WIDTH-1:0] rob_tag_in,
	input logic [STQ_SIZE-1:0] store_mask,

	// signals to store addresses from an AGU
	input logic agu_address_valid,
	input logic [XLEN-1:0] agu_address_data,
	input logic [ROB_TAG_WIDTH-1:0] agu_address_rob_tag,	// use to identify which

	// signals to indicate a load has been fired
	input logic load_executed,
	input logic [ROB_TAG_WIDTH-1:0] load_executed_rob_tag,

	// signals from the memory interface to designate a succeeded load
	// the load_succeeded_rob_tag is tracked by cache miss registers in
	// the caches
	input logic load_succeeded,				// bool to say if a load succeeded
	input logic [ROB_TAG_WIDTH-1:0] load_succeeded_rob_tag,	// ROB tag of the succeeded load

	// rob signals to know when loads commit
	input logic rob_commit,
	input logic [ROB_TAG_WIDTH-1:0] rob_commit_tag,

	// each bit determines if that entry experienced an order failure
	// multiple loads may have their order failures set at once, if they
	// all loaded before the committing store
	input logic [LDQ_SIZE-1:0] order_failures,

	// circular buffer pointers
	output load_queue_entry [LDQ_SIZE-1:0] load_queue_entries,
	output logic [$clog2(LDQ_SIZE)-1:0] head,
	output logic [$clog2(LDQ_SIZE)-1:0] tail,

	output logic full
	// TODO flush signals
	);

	// loop iterator
	integer i;

	always_ff @ (posedge clk) begin
		if (!reset) begin
			head <= 0;
			tail <= 0;

			for (i = 0; i < LDQ_SIZE; i = i + 1) begin
				clear_entry(i);
			end
		end else begin
			// place a new load instruction in the load buffer
			if (alloc_ldq_entry) begin
				load_queue_entries[tail].valid <= 1;
				load_queue_entries[tail].rob_tag <= rob_tag_in;
				load_queue_entries[tail].store_mask <= store_mask;
				tail <= tail + 1;
			end

			// if the entry at the head is committed, free it and increment head
			if (load_queue_entries[head].committed) begin
				clear_entry(int'(head));
				head <= head + 1;
			end

			// TODO:
			// - order_fail
			//	- "To discover ordering failures, when a store
			//	commits, it checks the entire LDQ for any
			//	address matches. If there is a match, the
			//	store checks to see if the load has executed,
			//	and if it got its data from memory or if the
			//	data was forwarded from an older store. In
			//	either case, a memory ordering failure has
			//	occurred."
			//	- needs to be able to update all or multiple
			//	entries in one cycle
			// - forward_stq_data
			// - forward_stq_index

			// loop to do operations on every entry
			for (i = 0; i < LDQ_SIZE; i = i + 1) begin	// each entry in the buffer makes this comparison
				// READ ADDRESS FROM THE AGU
				// if the address from the AGU is to be read and the ROB tag matches
				if (load_queue_entries[i].valid && agu_address_valid && agu_address_rob_tag == load_queue_entries[i].rob_tag) begin
					// if match, update address and declare it to be valid
					load_queue_entries[i].address <= agu_address_data;
					load_queue_entries[i].address_valid <= 1;
				end

				if (load_queue_entries[i].valid && load_executed && load_executed_rob_tag == load_queue_entries[i].rob_tag) begin
					load_queue_entries[i].executed <= 1;
				end

				if (load_queue_entries[i].valid && load_succeeded && load_succeeded_rob_tag == load_queue_entries[i].rob_tag) begin
					load_queue_entries[i].succeeded <= 1;
				end

				/*
				* here is a potential flaw of my design: I track that this
				* load has been committed this cycle so that the queue entry
				* can be freed the next cycle at the earliest.  One could
				* assume that the commit coming from the ROB is guaranteed to
				* be the load at the head of the queue.  But since I haven't
				* defined hardware to check that, I'm not making that
				* assumption.  Instead, I'm just going to have the head check
				* that it's pointing to a committed entry before clearing the
				* entry and incrementing.
				*/
				if (load_queue_entries[i].valid
						&& rob_commit
						&& rob_commit_tag == load_queue_entries[i].rob_tag) begin
					load_queue_entries[i].committed <= 1;
				end

				// set the order fail bit of this entry if it was detected by the searcher
				load_queue_entries[i].order_fail <= load_queue_entries[i].order_fail | order_failures[i];
			end
		end
	end

	// Since the tail pointer points to the next available entry in the
	// buffer, if that entry has the valid bit set, there are no more
	// available entries and the buffer is full.
	assign full = load_queue_entries[tail].valid;

	function void clear_entry(integer index);
		load_queue_entries[index].valid <= 0;
		load_queue_entries[index].address <= 0;
		load_queue_entries[index].address_valid <= 0;
		load_queue_entries[index].executed <= 0;
		load_queue_entries[index].succeeded <= 0;
		load_queue_entries[index].committed <= 0;
		load_queue_entries[index].order_fail <= 0;
		load_queue_entries[index].store_mask <= 0;
		load_queue_entries[index].forward_stq_data <= 0;
		load_queue_entries[index].forward_stq_index <= 0;
		load_queue_entries[index].rob_tag <= 0;
	endfunction
endmodule
